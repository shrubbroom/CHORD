`include "pipeline.v"
`include "interface_input.v"
module top();
   /*dummy top*/
endmodule // top
